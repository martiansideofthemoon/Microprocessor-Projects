library std;
library ieee;
use ieee.std_logic_1164.all;
package CacheComponent is

type CacheArray is array(0 to 15) of std_logic_vector(32 downto 0);

constant INIT_CACHE : CacheArray := (
  0 => "000000000000000000000000000000000",
  1 => "000000000000000000000000000000000",
  2 => "000000000000000000000000000000000",
  3 => "000000000000000000000000000000000",
  4 => "000000000000000000000000000000000",
  5 => "000000000000000000000000000000000",
  6 => "000000000000000000000000000000000",
  7 => "000000000000000000000000000000000",
  8 => "000000000000000000000000000000000",
  9 => "000000000000000000000000000000000",
  10 => "000000000000000000000000000000000",
  11 => "000000000000000000000000000000000",
  12 => "000000000000000000000000000000000",
  13 => "000000000000000000000000000000000",
  14 => "000000000000000000000000000000000",
  15 => "000000000000000000000000000000000"
);

end CacheComponent;
