
library ieee;
use ieee.std_logic_1164.all;
library work;
use work.ProcessorComponents.all;
entity ResetMemory is
  port (
    memory: out MemArray
  );
end entity ResetMemory;

architecture Struct of ResetMemory is
begin
  memory(0) <= "00011110";
  memory(1) <= "00010010";
  memory(2) <= "00111110";
  memory(3) <= "01100000";
  memory(4) <= "11101000";
  memory(5) <= "00001000";
  memory(6) <= "01000010";
  memory(7) <= "00000010";
  memory(8) <= "10100000";
  memory(9) <= "00000110";
  memory(10) <= "01011000";
  memory(11) <= "00000100";
  memory(12) <= "00111110";
  memory(13) <= "01110000";
  memory(14) <= "11000000";
  memory(15) <= "00011101";
  memory(16) <= "10011101";
  memory(17) <= "01000001";
  memory(18) <= "00001000";
  memory(19) <= "00000000";
  memory(20) <= "10001010";
  memory(21) <= "00001101";
  memory(22) <= "00001001";
  memory(23) <= "00000000";
  memory(24) <= "00001010";
  memory(25) <= "00100000";
  memory(26) <= "10001000";
  memory(27) <= "00001101";
  memory(28) <= "00001001";
  memory(29) <= "00100000";
  memory(30) <= "11111111";
  memory(31) <= "00110000";
  memory(32) <= "10011110";
  memory(33) <= "01010001";
  memory(34) <= "10001000";
  memory(35) <= "00001101";
  memory(36) <= "10000010";
  memory(37) <= "11000011";
  memory(38) <= "00001000";
  memory(39) <= "00001011";
  memory(40) <= "00000010";
  memory(41) <= "10000000";
  memory(42) <= "00001000";
  memory(43) <= "00001011";
  memory(44) <= "10000000";
  memory(45) <= "10010001";
  memory(46) <= "00000000";
  memory(47) <= "00000000";
  memory(48) <= "00000000";
  memory(49) <= "00000000";
  memory(50) <= "00000000";
  memory(51) <= "00000000";
  memory(52) <= "00000000";
  memory(53) <= "00000000";
  memory(54) <= "00000000";
  memory(55) <= "00000000";
  memory(56) <= "00000000";
  memory(57) <= "00000000";
  memory(58) <= "00000000";
  memory(59) <= "00000000";
  memory(60) <= "00000000";
  memory(61) <= "00000000";
  memory(62) <= "00000000";
  memory(63) <= "00000000";
  memory(64) <= "00000000";
  memory(65) <= "00000000";
  memory(66) <= "00000000";
  memory(67) <= "00000000";
  memory(68) <= "00000000";
  memory(69) <= "00000000";
  memory(70) <= "00000000";
  memory(71) <= "00000000";
  memory(72) <= "00000000";
  memory(73) <= "00000000";
  memory(74) <= "00000000";
  memory(75) <= "00000000";
  memory(76) <= "00000000";
  memory(77) <= "00000000";
  memory(78) <= "00000000";
  memory(79) <= "00000000";
  memory(80) <= "00000000";
  memory(81) <= "00000000";
  memory(82) <= "00000000";
  memory(83) <= "00000000";
  memory(84) <= "00000000";
  memory(85) <= "00000000";
  memory(86) <= "00000000";
  memory(87) <= "00000000";
  memory(88) <= "00000000";
  memory(89) <= "00000000";
  memory(90) <= "00000000";
  memory(91) <= "00000000";
  memory(92) <= "00000000";
  memory(93) <= "00000000";
  memory(94) <= "00000000";
  memory(95) <= "00000000";
  memory(96) <= "00000000";
  memory(97) <= "00000000";
  memory(98) <= "00000000";
  memory(99) <= "00000000";
  memory(100) <= "00000000";
  memory(101) <= "00000000";
  memory(102) <= "00000000";
  memory(103) <= "00000000";
  memory(104) <= "00000000";
  memory(105) <= "00000000";
  memory(106) <= "00000000";
  memory(107) <= "00000000";
  memory(108) <= "00000000";
  memory(109) <= "00000000";
  memory(110) <= "00000000";
  memory(111) <= "00000000";
  memory(112) <= "00000000";
  memory(113) <= "00000000";
  memory(114) <= "00000000";
  memory(115) <= "00000000";
  memory(116) <= "00000000";
  memory(117) <= "00000000";
  memory(118) <= "00000000";
  memory(119) <= "00000000";
  memory(120) <= "00000000";
  memory(121) <= "00000000";
  memory(122) <= "00000000";
  memory(123) <= "00000000";
  memory(124) <= "00000000";
  memory(125) <= "00000000";
  memory(126) <= "00000000";
  memory(127) <= "00000000";
end Struct;